module vit
